module Adder_PC
(
	data1_i,	// program counter now
	data2_i,	// 4
	data_o
);

input	[31:0]		data1_i;
input	[31:0]		data2_i;
output	[31:0]		data_o;

assign	data_o		= data1_i + data2_i;

endmodule